module Cfu (
    input               cmd_valid,
    output           cmd_ready,
    input      [9:0]    cmd_payload_function_id,
    input      [31:0]   cmd_payload_inputs_0,
    input      [31:0]   cmd_payload_inputs_1,
    output reg          rsp_valid,
    input               rsp_ready,
    output reg [31:0]   rsp_payload_outputs_0,
    input               reset,
    input               clk
);

    // reg [8:0] InputOffset = $signed(9'd128), FilterOffset = $signed(9'd0);
    localparam InputOffset = $signed(9'd128);

    // SIMD multiply step:
    wire signed [15:0] prod_0, prod_1, prod_2, prod_3;
    // wire signed [8:0] cur_offset;

    // assign cur_offset = |cmd_payload_inputs_0[31:8]?InputOffset:FilterOffset;

    assign prod_0 = ($signed(cmd_payload_inputs_0[7 : 0]) + InputOffset)
                  * $signed(cmd_payload_inputs_1[7 : 0]);
    assign prod_1 = ($signed(cmd_payload_inputs_0[15 : 8]) + InputOffset)
                  * $signed(cmd_payload_inputs_1[15 : 8]);
    assign prod_2 = ($signed(cmd_payload_inputs_0[23 : 16]) + InputOffset)
                  * $signed(cmd_payload_inputs_1[23 : 16]);
    assign prod_3 = ($signed(cmd_payload_inputs_0[31 : 24]) + InputOffset)
                  * $signed(cmd_payload_inputs_1[31 : 24]);

    wire signed [31:0] sum_prods;
    assign sum_prods = prod_0 + prod_1 + prod_2 + prod_3;

    // Only not ready for a command when we have a response.
    assign cmd_ready = ~rsp_valid;

    always @(posedge clk) begin
        if (reset) begin
          rsp_payload_outputs_0 <= 32'b0;
          rsp_valid <= 1'b0;
        end else if (rsp_valid) begin
          rsp_valid <= ~rsp_ready;
        end else if(cmd_valid) begin
          rsp_valid <= 1'b1;
          rsp_payload_outputs_0 <= |cmd_payload_function_id[9:3]
          ? 32'b0
          : rsp_payload_outputs_0 + sum_prods;
        end
    end
endmodule